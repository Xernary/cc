    Mac OS X            	   2   �      �                                      ATTR       �   �   *                  �     com.apple.lastuseddate#PS       �     com.dropbox.attrs    ��5b    "�[,    

B��J�     ����ӹ