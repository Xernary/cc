    Mac OS X            	   2       F                                      ATTR      F   �   f                  �     com.apple.lastuseddate#PS       �   <  com.apple.quarantine   ,     com.dropbox.attrs    ��|b    ��    q/0081;627cc332;Chrome;90BD033F-86EE-4ECF-8155-39D75D8C4040 

B��J�     ������